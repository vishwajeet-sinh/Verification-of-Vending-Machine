package vend_pkg;

import uvm_pkg::*;
`include "trans.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "monitor_dut.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"

endpackage
